
module ALTCLKCTRL (
	inclk,
	outclk);	

	input		inclk;
	output		outclk;
endmodule
