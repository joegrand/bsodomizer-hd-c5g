
module sfl (
	noe_in);	

	input		noe_in;
endmodule
